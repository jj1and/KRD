`ifndef __FEE_CONFIG_VH__
`define __FEE_CONFIG_VH__

// Trigger parameters
`define ADC_RESOLUTION_WIDTH 12
`define SAMPLE_WIDTH 16

`endif