`timescale 1 ns / 1ps

module SFP_module_IF # (

)
(

);

endmodule